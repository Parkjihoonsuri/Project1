module stop_watch_top(
    input clk,
    input reset_p,
    input [1:0] btn,
    output [3:0] com,
    output [7:0] seg_7,
    output [7:0] led_bar
    );
    
    reg[25:0] clk_div;
    wire btn_start, start_stop;
    wire [1:0] debounced_btn;
    always @(posedge clk) clk_div <= clk_div + 1;

    d_flip_flop_p dff0(.d(btn[0]), .clk(clk_div[16]), .reset_p(reset_p), .q(debounced_btn[0]));
    edge_detector_n ed_start(.clk(clk), .cp_in(debounced_btn[0]), .reset_p(reset_p), .p_edge(btn_start));
    t_flip_flop_p (.clk(clk), .t(btn_start), .reset_p(reset_p), .q(start_stop));
    
    wire lap, btn_lap;
    d_flip_flop_p dff1(.d(btn[1]), .clk(clk_div[16]), .reset_p(reset_p), .q(debounced_btn[1]));
    edge_detector_n ed_lap(.clk(clk), .cp_in(debounced_btn[1]), .reset_p(reset_p), .p_edge(btn_lap));
    t_flip_flop_p (.clk(clk), .t(btn_lap), .reset_p(reset_p), .q(lap));
    
    assign led_bar[0] = debounced_btn[1];
    assign led_bar[1] = btn_lap;
    assign led_bar[2] = lap;
    
    wire clk_usec;
    clock_usec usec_clk(.clk(clk), .reset_p(reset_p), .clk_usec(clk_usec));
    wire clk_msec;
    clock_msec msec_clk(.clk(clk), .reset_p(reset_p), .clk_usec(clk_usec), .clk_msec(clk_msec));
    wire clk_sec;
    
    wire clk_start;
    assign clk_start = start_stop ? clk_msec : 1'b0; // ����/���� ��ư���� msec Ŭ�� ����

    clock_sec sec_clk(.clk(clk), .reset_p(reset_p), .clk_msec(clk_start), .clk_sec(clk_sec));
    wire clk_min;
    clock_min min_clk(.clk(clk), .clk_sec(clk_sec), .reset_p(reset_p), .clk_min(clk_min));
    
    wire [3:0] sec1, sec10, min1, min10;

    counter_dec_60(.clk(clk), .reset_p(reset_p), .clk_time(clk_sec), .dec1(sec1), .dec10(sec10));
    counter_dec_60(.clk(clk), .reset_p(reset_p), .clk_time(clk_min), .dec1(min1), .dec10(min10));

    reg [15:0] lap_value;
    always @(posedge clk or posedge reset_p) begin
        if (reset_p) lap_value <= 0;
        else if (btn_lap) lap_value <= {sec10, sec1, min10, min1}; // ���÷��� ���� �ʿ� �и��ʷ� ������Ʈ
    end

    wire [15:0] value;
    assign value = lap ? lap_value : {sec10, sec1, min10, min1}; // ���÷��� ���� �ʿ� �и��ʷ� ǥ��

    fnd_4digit_cntr fnd_cntr(.clk(clk), .reset_p(reset_p), .value(value), .com(com), .seg_7(seg_7));

    // ������ ������ ��� �ν��Ͻ�ȭ �κ� (���� �� ��Ʈ ������ ���� ���� ��ġ�ϰ� ���� �ʿ�)

endmodule
